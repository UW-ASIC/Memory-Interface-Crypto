module spi_controller (
    input wire clk, 
    input wire rst_n,
    input wire done,
    input wire [7:0] address, //or [23:0] address
    input wire [7:0] data
);
    
endmodule